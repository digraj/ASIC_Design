// $Id: $
// File name:   flex_stp_sr.sv
// Created:     1/26/2017
// Author:      Kunwar Digraj Singh Jain
// Lab Section: 5
// Version:     1.0  Initial Design Entry
// Description: serial to parallel shift register

module flex_stp_sr 
#(
	parameter 	NUM_BITS = 4,
			SHIFT_MSB = 1 
)
(
	input wire 	clk,
			n_rst,
			shift_enable,
			serial_in, 
	output reg	[NUM_BITS-1:0] parallel_out,
	output reg 	byte_rcv
);

	reg [NUM_BITS-1:0]mid_output ;
	
	always_comb
	begin
		if (!shift_enable == 1'b0)
		begin
			mid_output = parallel_out ;
		end
		else if (!shift_enable == 1'b1)
		begin
			if (SHIFT_MSB == 1'b1) 
			begin
				mid_output = {parallel_out[NUM_BITS-2:0], serial_in} ;
			end
			else 
			begin
				mid_output = {serial_in, parallel_out[NUM_BITS-1:1]} ;
			end		
		end
	end

	always_ff @ (posedge clk, negedge n_rst)
	begin
		if (n_rst == 1'b0)
		begin
			byte_rcv = 0 ;
			parallel_out <= '1 ;	
		end
		else 
		begin
			byte_rcv <= shift_enable ;
			parallel_out <= mid_output ;
		end
	end

endmodule
